package macGenClassPckg;
	`include "macGenClass.sv";
endpackage
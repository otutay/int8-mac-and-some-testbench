package im2ColGenClassPckg;
	`include "im2ColGenClass.sv";
endpackage
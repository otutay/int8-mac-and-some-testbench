otutay@eotPc.6968:1576782802
package macMonitorClassPckg;
	`include "macMonitorClass.sv";
endpackage
package macTestEnvClassPckg;
	`include "macTestEnvClass.sv";
endpackage
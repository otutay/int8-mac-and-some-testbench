package generatorPckg;
	`include "generator.sv";
endpackage
otutay@eotPc.9302:1576782802
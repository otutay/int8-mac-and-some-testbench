package macTransClassPckg;
	`include "macTransClass.sv";
endpackage
package environmentPckg;
	`include "environment.sv";
endpackage
package macScoreClassPckg;
	`include "macScoreClass.sv";
endpackage
package transactionPckg;
	`include "transaction.sv";
endpackage : transactionPckg
package macDriverClassPckg;
	`include "macDriverClass.sv";
endpackage
package driverPckg;
	`include "driver.sv";
endpackage
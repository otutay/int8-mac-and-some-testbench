package tilePckg;
	parameter cNumOfRam = 32;
	parameter cNumOfMul = 12;

endpackage
import macPckg::*;

class macTransClass;
	rand tMultIn iData;
	tMultOut oData;

	// no constraint as it accept every range of inputs.
	// constraint dvAllZero { iData.dv == 1'b0;
		
	// }
endclass : macTransClass
package im2ColTransClassPckg;
	`include "im2ColTransClass.sv";
endpackage
package im2ColDrivClassPckg;
	`include "im2ColDrivClass.sv";
endpackage
package im2ColEnvClassPckg;
	`include "im2ColEnvClass.sv";
endpackage